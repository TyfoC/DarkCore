LEF0 �    @ 0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     6          0        "  |       (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �*  �   ����U�����hG"@ ��  ���  @ ��Ph`"@ ��  ��� @ ��Ph�"@ ��  ��� @ ��Ph�"@ �  ��� @ ��Ph�"@ �  ��� @ ��Ph�"@ �  ��� @ ��Ph�"@ �i  ��� @ ��Ph�"@ �S  ��� @ ��Ph#@ �=  ���  @ ��Ph4#@ �'  ���$ @ ��Ph`#@ �  ���( @ ��Ph�#@ ��  ���, @ ��Ph�#@ ��  ����ÍL$����q�U��WSQ��  ��jj h�#@ �  ����h$@ �  ����h�  h (@ ��  ���  @ ��j Ph (@ �s  ��������t�j���볡 @ ��j Ph (@ �K  ��������t(��  ��j j ��  ����j j��  ���j���� @ ��j Ph (@ �  ����������   �E�    ��E�E� (@ � < t!�E� (@ � <	t�E� (@ � ��u���E�E� (@ � < t�E� (@ � <	u�E� (@ � ��uӋE� (@ ��P�n  ����h
$@ �^  ������� @ ��j Ph (@ �O  ��������tj��h    ��  ���E��}� t�$@ ��$@ ��Ph$@ �  �����u��f  ����t�$@ ��$@ ��Ph+$@ ��  ���,���� @ ��j Ph (@ ��  ��������t
��  ����� @ ��j Ph (@ �  ��������t
�  ������ @ ��j Ph (@ �n  ��������t8��  �E����u�h>$@ �R  ���}� ��������u��#  ���}���� @ ��j Ph (@ �  ����������   �E�    ��E��E� (@ � < t!�E� (@ � <	t�E� (@ � ��u���E��E� (@ � < t�E� (@ � <	u�E� (@ � ��uӋE� (@ � ��������E� (@ ��P�E  �������������hT$@ �j  �������  @ ��j Ph (@ �E  ����������  �  �Eč�k����   �    �߉�����k���P�u���  ������t��h|$@ ��  ���  �������)  � �߉���Z  ��������P�  ���E���u�E��U���Ph�$@ �  ���7�E�<u�E��U���Ph�$@ �  ����E�<u��h�$@ �Z  ���E��U�	Ѕ���   ��h�$@ �:  ���E��U�����`���ǅd���    ��`�����d���	Ѕ�t��h�$@ ��  ���E��U�����X���ǅ\���    ��X�����\���	Ѕ�t��h�$@ ��  ���E��U�����P���ǅT���    ��P�����T���	Ѕ�t��h�$@ �  ����h%@ �y  ����h
$@ �i  ����������P��k���P�p  ����������}� ��������u��/  �������$ @ ��j Ph (@ �!
  ����������  �E�    ��E܋E� (@ � < t!�E� (@ � <	t�E� (@ � ��u���E܋E� (@ � < t�E� (@ � <	u�E� (@ � ��uӋE� (@ � ��������E܍� (@ ��������RP�  ������������  ��������Ph%@ �d  ���E���u�%@ ��%@ ��Ph#%@ �@  ���E��U�	Ѕ���   ��h.%@ �   ����h�$@ ��  ���E��U�����H���ǅL���    ��H�����L���	Ѕ�t��h�$@ �  ���E��U�����@���ǅD���    ��@�����D���	Ѕ�t��h�$@ �  ���E��U�����8���ǅ<���    ��8�����<���	Ѕ�t��h�$@ �I  ����h%@ �9  ����h
$@ �)  ���E���u�E��U���RPh;%@ �   ����E��U���RPhL%@ �  ���U��E���RPhh%@ ��  ���U��E���RPh�%@ ��  ���U��E���RPh�%@ �  ����E� (@ ��Ph�%@ �  ����h)  j ������P�R  ��������( @ ��j Ph (@ �e  ���������  �E�    ��E؋E� (@ � < t!�E� (@ � <	t�E� (@ � ��u���E؋E� (@ � < t�E� (@ � <	u�E� (@ � ��uӋE� (@ � ���1����E؍� (@ ���E�PR�$  ���Eȃ}� u��h &@ �  ��������E�    ��UȋE�Њ ����P�\  ���EԋE�9E�r܃}� t���u��Z  ����h
$@ �K  �������, @ ��j Ph (@ �<  ����������   �E�    ��EЋE� (@ � < t!�E� (@ � <	t�E� (@ � ��u���EЋE� (@ � < t�E� (@ � <	u�E� (@ � ��uӋE� (@ � �������EЍ� (@ ���E�PR��  ���Ẽ}� u��h &@ �  ��������E���j
P�u��  ���}� t���u��J  ����h
$@ �;  ������� (@ ��������  @ ��Ph (@ h &@ �$  ���g���U��� �E�    �E����t
�E����u@�E�E�E�E��%�E���    �E�ЋU���    �U�ʋ ��E��E��9E�r���E����t
�E����u<�E�E��E�E��"�E���E��E���E��f�f��E��E��9E�r��.�E�E��E�E���U�E�ЋM��U�ʊ ��E��E�;Erᐐ��U���$�E�E��E�    �E����t
�E����uN�E�E��U܉���������E���	��E�	ЉE���E���    �E�E��E��E��9E�r��o�E����t
�E����u9�E�E��U܉����f�E���E���E��f�E�f��E��E��9E�r��!�E�E���U��E�E܈�E��E�;Er萐��U��� �E�    �E����t
�E����uN�E�E�E�E��0�E���    �E�Ћ�E���    �E�ȋ 9�t� �   �E��E��9E�r��   �E����t
�E����uD�E�E��E�E��*�E���E��f��E�����E��f� f9�t� �F�E��E��9E�r��5�E�E��E�E���U��E�Њ�M�E�Ȋ 8�t� ��E��E�;Erٰ��U����}w������(�E�   ��E��E�    �u�E�} ����u�E��ÐU����E��y�؉E��u�u���������U����}v�}v� �   �} u�E� 0�E@�  ��r�E�E��E�   ��E��E��    �u�E��}� ����u�U�E�ЉE�E��  �M��)�E�    �u�Њ�l&@ �E��E�    �u�E�M�} uѰ��U��} y�E� -�]�E�E�uP�u�8������ÐU����E�    �6�U�E�Њ <`~%�U�E�Њ <z�U�E�Њ�M�E�ȃ�_��E��U�E�Њ ��u����ÐU����E�    �6�U�E�Њ <@~%�U�E�Њ <Z�U�E�Њ�M�E�ȃ� ��E��U�E�Њ ��u����ÐU����E�    ��E��U�E�Њ ��u�E��ÐU����E�    �U�E�Њ�M�E�Ȋ 8�t� ��U�E�Њ ��t�E��ѐ��ÐU����u�������E��u�|������E��U�E��9E�r�}�u������d�E�)E��O�E��E�    �&�U�E�EЊ�M�E�Ȋ 8�t�E� ��E��U�E�Њ ��ù}� t�E��E�E9E�s��������U����u��������E�E;E�r� �N�} u�E�+E�E��U�E�9E�s	�E�+E�E�U�EЃ��uP�u��������U�E��  ���U�� 0@ ��v������^� 0@ �������� *@ �E�� 0@ ��������*@ �E�� 0@ ��������*@ �E�� 0@ @� 0@ �    ]�U���� 0@ �E�} ��   �F�U������ *@ � ��t/�U������ *@ ��M������*@ � ��P�҃��E�P��U������u��p�U������ *@ � 9EuF�U������ *@ ��M������*@ � ��P�҃��U������ *@ �     �E�P��U������u���U��E� ������]�U��E� �]�U��]�U��E�    �u�ЋU)E�]�U����E�    �u�U��E�)E�E;Es	�E    ��E)E�E��U���(���u�=  ���E�    �E�    �E�    �8  �E�U�E�Њ <t*�U�E�Њ <
t�U�E�Њ < t�U�E�Њ <	u�E�;Er��E�;E��  �E�E���E��U�E�Њ < t2�U�E�Њ <	t$�U�E�Њ <t�U�E�Њ <
t�E�;Er��E�+E�E�E�@��P��  ���E��U�E�E����u�RP�������U��E���  �E�@�E�E�;E�Z  ��E�U�E�Њ <t*�U�E�Њ <
t�U�E�Њ < t�U�E�Њ <	u�E�;Er��E�;E�  �U�E�Њ <=u�E���E�U�E�Њ <t*�U�E�Њ <
t�U�E�Њ < t�U�E�Њ <	u�E�;Er��E�9E��   �E�E���E��U�E�Њ <t�U�E�Њ <
t�E�;ErًE�+E�E�E��P��  ���E�U�E�E���u�RP��������U�E���  ���E�P�u�Y  ���E�@�E��E�    �E�E��E�;E������
���������E�� U������u��  ���E��E�    �   ���u��u��  ��� ������t#���u��u��  ��� ��t��P�*  �����u��u�  ���@������t$���u��u�  ���@��t��P��  ���E�E�;E��q�������U��    �    ����]�U��    �   ����]�U����   �    �U��E��E��ÐU����   �   �U��E��}����ÐU��   �    ����]�U����   �   �U��E��E��ÐU��S�   �   �U�]�쐋]���U����E�E��   �   �U�����U��   �   �U��]ÐU��U�   �   ��]ÐU��VS�   �   �U�]�u��[^]ÐU��S�   �    �U�]�쐋]���U��   �   ����]�U����   �    ����E�E��P�������E��E�@��P�  ���E�E��P�E��RP�u��,������E���U����   �   �U��E��}����ÐU��S���]�   �   �U��E��}����]���U��S���U�]�   �   ��E��}����]���U��S�]�   �   �U�쐋E�]��� �U����U�   �   ��ʉE��U��E�U���E���U����   �    ����E��E���U����   �    �U��E��E���U����   �    �U��E��E���U��   �   �U��]�U��   �   �U��]�U��   �   �U��]�U��   �   �U��]�U����E�     �E�@    �E�@    ��jP�b������E��E� ��t�E�@
   �E�@    ���� U��S���E� ��u� ��   �E�P�E�@9���   �E�@��
=���w����������P��������E�}� u� �|�E�@�P
�E�P�E�@��    �E� ��RP�u���������E� ��t�E� ��P��������E�U��E��E�@�H�U�J����E�P� ��Q��]��� U��E�@]� U��E� �U���]�                                                                                                                   "@ "@ "@ "@ "@  "@ '"@ ,"@ /"@ 2"@ 7"@ ?"@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 help clear echo vmtest shutdown reboot path cd ls info txtread hexread Supported commands:
    	%s - get info about commands
 	%s - clear terminal
 	%s <text> - echo some text
    	%s - test VMM memory allocation
 	%s - shutdown
 	%s - reboot
 	%s - get current path
 	%s <path> - set current path
 	%s - show objects in current directory
   	%s <path> - show file system object information
  	%s <path> - show txt file content
    	%s <path> - show hex file content
    Welcome to DarkCore Shell v%u.%u
 #  
 yes no Memory allocated: %s
 Memory freed: %s
 Current path: `%s`
  %a0CError: invalid directory path!
    Error: cannot create directory iterator!
  - file (%u bytes)  - directory (%u elements)  - symbolic link  [ SYSTEM  READ_ONLY  HIDDEN  ] Name: `%s`
 file directory Type: %s
 Attributes:  Size: %u bytes
 Files & Folders Count: %u
 Creation Date & Time: %x %x
   Last Read Date & Time: %x %x
  Last Write Date & Time: %x %x
 %a0CError: cannot get information about %a0E`%s`%a0C!
 %a0CError: cannot read file!
  %a0CError: unknown command: `%s` %a07(Type `%a0A%s`%a07 to get info)%a0C!
 0123456789ABCDEF